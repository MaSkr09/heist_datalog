----------------------------------------------------------------------------------
-- MIT License
-- 
-- Copyright (c) 2022 Martin Skriver
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
----------------------------------------------------------------------------------
-- Company: University of Southern Denmark
-- Engineer: Martin Skriver
-- Contact: maskr@mmmi.sdu.dk
--
-- Description: 
-- BRAM instantiation for HEIST
--
----------------------------------------------------------------------------------

--------------------------------------------------------------------------
-- DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width --
-- ===============|===========|===========|===============|=============--
--          19-36 |    "36Kb" |      1024 |        10-bit |       4-bit --
--          10-18 |    "36Kb" |      2048 |        11-bit |       2-bit --
--          10-18 |    "18Kb" |      1024 |        10-bit |       2-bit --
--            5-9 |    "36Kb" |      4096 |        12-bit |       1-bit --
--            5-9 |    "18Kb" |      2048 |        11-bit |       1-bit --
--            3-4 |    "36Kb" |      8192 |        13-bit |       1-bit --
--            3-4 |    "18Kb" |      4096 |        12-bit |       1-bit --
--              2 |    "36Kb" |     16384 |        14-bit |       1-bit --
--              2 |    "18Kb" |      8192 |        13-bit |       1-bit --
--              1 |    "36Kb" |     32768 |        15-bit |       1-bit --
--              1 |    "18Kb" |     16384 |        14-bit |       1-bit --
--------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------
-- Libraries 
-----------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VComponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

-----------------------------------------------------------------------------------------------------
-- Ports and generics
-----------------------------------------------------------------------------------------------------
entity true_dual_port_bram_inst is
    generic (
        mem_size            : string := "36Kb"; -- Target BRAM, "18Kb" or "36Kb"
        read_width_a        : integer := 8;     -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        read_width_b        : integer := 8;     -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        write_width_a       : integer := 8;     -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        write_width_b       : integer := 8;     -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        addr_width_a        : integer := 12;    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        addr_width_b        : integer := 12;    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        write_en_width_a    : integer := 1;     -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        write_en_width_b    : integer := 1      -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
    );
    Port ( 
        CLKA_in             : in STD_LOGIC;           -- 1-bit input port-A clock
        DOA_out             : out STD_LOGIC_VECTOR((read_width_a-1) downto 0);      -- Output port-A data, width defined by READ_WIDTH_A parameter
        ADDRA_in            : in STD_LOGIC_VECTOR((addr_width_a-1) downto 0);       -- Input port-A address, width defined by Port A depth
        DIA_in              : in STD_LOGIC_VECTOR((write_width_a-1) downto 0);                 -- Input port-A data, width defined by WRITE_WIDTH_A parameter
        ENA_in              : in STD_LOGIC;                                         -- 1-bit input port-A enable
--        REGCEA_in           : in STD_LOGIC;                                         -- 1-bit input port-A output register enable
        RSTA_in             : in STD_LOGIC;                                         -- 1-bit input port-A reset
        WEA_in              : in STD_LOGIC_VECTOR((write_en_width_a-1) downto 0);   -- Input port-A write enable, width defined by Port A depth

        CLKB_in             : in STD_LOGIC;           -- 1-bit input port-B clock
        DOB_out             : out STD_LOGIC_VECTOR((read_width_b-1) downto 0);      -- Output port-B data, width defined by READ_WIDTH_B parameter
        ADDRB_in            : in STD_LOGIC_VECTOR((addr_width_b-1) downto 0);       -- Input port-B address, width defined by Port B depth
        DIB_in              : in STD_LOGIC_VECTOR((write_width_b-1) downto 0);                 -- Input port-B data, width defined by WRITE_WIDTH_B parameter
        ENB_in              : in STD_LOGIC;                                         -- 1-bit input port-B enable
--        REGCEB_in           : in STD_LOGIC;                                         -- 1-bit input port-B output register enable
        RSTB_in             : in STD_LOGIC;                                         -- 1-bit input port-B reset
        WEB_in              : in STD_LOGIC_VECTOR((write_en_width_b-1) downto 0)    -- Input port-B write enable, width defined by Port B depth

    );
end true_dual_port_bram_inst;

architecture Behavioral of true_dual_port_bram_inst is

begin
BRAM_TDP_MACRO_inst : BRAM_TDP_MACRO
    generic map (
        BRAM_SIZE           => mem_size,        -- Target BRAM, "18Kb" or "36Kb"
        DEVICE              => "7SERIES",       -- Target Device: "VIRTEX5", "VIRTEX6", "7SERIES", "SPARTAN6"
        DOA_REG             => 0,               -- Optional port A output register (0 or 1)
        DOB_REG             => 0,               -- Optional port B output register (0 or 1)
        INIT_A              => X"000000000",    -- Initial values on A output port
        INIT_B              => X"000000000",    -- Initial values on B output port
        INIT_FILE           => "NONE",
        READ_WIDTH_A        => read_width_a,    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH_B        => read_width_b,    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY",
        -- "GENERATE_X_ONLY" or "NONE"
        SRVAL_A             => X"000000000",    -- Set/Reset value for A port output
        SRVAL_B             => X"000000000",    -- Set/Reset value for B port output
        WRITE_MODE_A        => "WRITE_FIRST",   -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        WRITE_MODE_B        => "WRITE_FIRST",   -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        WRITE_WIDTH_A       => write_width_a,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        WRITE_WIDTH_B       => write_width_a,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        
        -- The following INIT_xx declarations specify the initial contents of the RAM
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",--X"1F1E1D1C1B1A191817161514131211100F0E0D0C0B0A09080706050403020100",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",--X"FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210FEDCBA9876543210",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",--X"505050504F4F4F4F4E4E4E4E4D4D4D4D4C4C4C4C4B4B4B4B4A4A4A4A49494949",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",--X"4848484847474747464646464545454544444444434343434242424241414141",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",--X"4848484847474747464646464545454544444444434343434242424241414141",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000", --8000000400000002800000040000000280000004000000028000000400000002
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000", 
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",--
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INIT_xx are valid when configured as 36Kb
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INITP_xx are for the parity bits
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INIT_xx are valid when configured as 36Kb
        INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
    )
    port map (
        DOA => DOA_out,             -- Output port-A data, width defined by READ_WIDTH_A parameter
        DOB => DOB_out,             -- Output port-B data, width defined by READ_WIDTH_B parameter
        ADDRA => ADDRA_in,         -- Input port-A address, width defined by Port A depth
        ADDRB => ADDRB_in,         -- Input port-B address, width defined by Port B depth
        CLKA => CLKA_in,           -- 1-bit input port-A clock
        CLKB => CLKB_in,           -- 1-bit input port-B clock
        DIA => DIA_in,             -- Input port-A data, width defined by WRITE_WIDTH_A parameter
        DIB => DIB_in,             -- Input port-B data, width defined by WRITE_WIDTH_B parameter
        ENA => ENA_in,             -- 1-bit input port-A enable
        ENB => ENB_in,             -- 1-bit input port-B enable
--        REGCEA => REGCEA_in,       -- 1-bit input port-A output register enable
--        REGCEB => REGCEB_in,       -- 1-bit input port-B output register enable
        REGCEA => '0',       -- 1-bit input port-A output register enable
        REGCEB => '0',       -- 1-bit input port-B output register enable
        RSTA => RSTA_in,           -- 1-bit input port-A reset
        RSTB => RSTB_in,           -- 1-bit input port-B reset
        WEA => WEA_in,             -- Input port-A write enable, width defined by Port A depth
        WEB => WEB_in              -- Input port-B write enable, width defined by Port B depth
    );

end Behavioral;
